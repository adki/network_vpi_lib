//----------------------------------------------------------------------------
// Copyright (c) 2014 by Ando Ki.
// All rights are reserved by Ando Ki.
//----------------------------------------------------------------------------
// top.v
//----------------------------------------------------------------------------
// VERSION: 2014.06.24.
//----------------------------------------------------------------------------
module top;
    initial begin
        $dumpfile("wave.vcd");
        $dumpvars(0);
        if (1) test_ethernet;
        if (1) test_udp_ip_ethernet;
        #10; $finish(2);
    end
    //------------------------------------------------------------------------
    `include "top_tasks_ethernet.v"
    `include "top_tasks_udp_ip_ethernet.v"
endmodule
//----------------------------------------------------------------------------
// Revision history:
//
// 2014.06.24: Started by Ando Ki (andoki@gmail.com)
//----------------------------------------------------------------------------
